-- Greg Stitt
-- University of Florida
-- EEL 5934/4930 Reconfigurable Computing
--
-- File: tb.vhd
--
-- Description: This file implements a simple testbench for the Fibonacci
-- calculator. Note that this entity uses std_logic_arith in order to
-- illustrate a different package. I highly recommend using numeric_std
-- instead.   
--
-- Comments: Ideally, the individual tests could be made into a procedure to
-- avoid copy and pasting.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;

entity gray_tb is
end gray_tb;

architecture behavior of gray_tb is

  component gray2
    port( clk      : in  std_logic;
          rst      : in  std_logic;
          output   : out std_logic_vector(3 downto 0));
  end component;

  --Inputs
  signal clk : std_logic                     := '0';
  signal rst : std_logic                     := '1';

  --Outputs
  signal output : std_logic_vector(3 downto 0);

begin

  uut : gray2
    port map(clk, rst, output);

  -- toggle clock
  clk <= not clk after 50 ns;

  -- process to test different inputs
  process
  begin

    -- reset circuit  
    rst <= '1';
    wait for 200 ns;
    rst <= '0';
    wait until clk'event and clk = '1';
    U_STATE : for i in 0 to 18 loop
        wait until clk'event and clk = '1';
    end loop ; -- U_STATE  
    wait;
  end process;

end;
